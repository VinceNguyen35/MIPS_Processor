----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/17/2020 07:46:29 PM
-- Design Name: 
-- Module Name: SignExtend - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SignExtend is
    port(   Din : in STD_LOGIC_VECTOR ( 15 downto 0 );
            Dout : out STD_LOGIC_VECTOR ( 31 downto 0 )
    );
end SignExtend;

architecture Behavioral of SignExtend is
begin
    Dout(15 downto 0) <= Din;
    Dout(31 downto 16) <= (31 downto 16 => Din(15));
end Behavioral;
